`ifndef V5_CALC_TEST_LIB_SV
 `define V5_CALC_TEST_LIB_SV
package calc_test_lib;
`include "uvm_macros.svh" // Include the UVM macros
   import uvm_pkg::*;      // import the UVM library
   import calc_agent_pkg::*;
   `include "v5_calc_test_simple.sv"
   endpackage
`endif;
